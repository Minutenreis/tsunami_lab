netcdf artificialtsunami_displ_1000 {
dimensions:
	x = 5 ;
	y = 3 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = 3,4,5,6,7 ;

 y = 1,2,3 ;

 z = 0,1,2,3,4,
  	5,6,7,8,9,
	10,11,12,13,14;
}
