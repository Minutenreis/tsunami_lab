netcdf artificialtsunami_displ_1000 {
dimensions:
	x = 10 ;
	y = 5 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = 0,1,2,3,4,5,6,7,8,9 ;

 y = 0,1,2,3,4 ;

 z = 0,1,2,3,4,5,6,7,8,9,
    10,11,12,13,14,15,16,17,18,19,
    20,21,22,23,24,25,26,27,28,29,
    30,31,32,33,34,35,36,37,38,39,
    40,41,42,43,44,45,46,47,48,49;
}
