netcdf artificialtsunami_displ_1000 {
dimensions:
	x = 10 ;
	y = 5 ;
variables:
	float x(x) ;
	float y(y) ;
	float z(y, x) ;

// global attributes:
		:Conventions = "COARDS" ;
data:

 x = 0,1,2,3,4,5,6,7,8,9 ;

 y = 0,1,2,3,4 ;

 z = -10,-10,-10,-10,-10,-10,-10,-10,-10,-10,
 -10,-10,-10,-10,-10,-10,-10,-10,-10,-10,
 -10,-10,-10,-10,-10,-10,-10,-10,-10,-10,
 -10,-10,-10,-10,-10,-10,-10,-10,-10,-10,
 -10,-10,-10,-10,-10,-10,-10,-10,-10,-10;
}
